module my_xor (
  output f,
  input a, b, c
);

// assign f to be the xor of a, b, c
xor(f, a, b, c);

endmodule
